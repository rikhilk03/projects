/* packet_valid is high untill header to payload data goes low for parity
parity_done is high when router recieves the parity
data_in to capture the address of the destination(2 bit)
soft_reset_0,1,2 and fifo_full signals from the synchronizer
low_pkt_valid is negation of the pkt_valid that is when it is high it means it received the packet(header to payload)
packets are not pending (transfered from source to destination). if it is low it indicates not completely transferred.
fifo_empty_0,1,2 signals from respective fifo's 
remaining all signals are generated by the FSM
**write_enb_reg signal is high for three states (load_data, load_after_full, Load_priority)
**rst_int_reg  is high for check_parity_error state
**busy signal is high for all except decode address, load_data and load_priority
Task t1 :- for small packet data )the states chandges from (decode_addr-> load_first_data:load_data-> Load_priority-> check_parity_error-> decode_addr)
*/
module router_fsm(input clk, rst, pkt_valid, parity_done, input [1:0] data_in, input soft_reset_0,
					soft_reset_1, soft_reset_2, fifo_full, low_pkt_valid, fifo_empty_0,
					fifo_empty_1, fifo_empty_2, output busy, detect_add, ld_state, laf_state,
					full_state, write_enb_reg, rst_int_reg, lfd_state);

parameter DECODE_ADDRESS = 3'b000, WAIT_TILL_EMPTY = 3'b001, LOAD_FIRST_DATA = 3'b010, LOAD_DATA = 3'b011, 
		  LOAD_PARITY = 3'b100,  CHECK_PARITY_ERROR = 3'b101, FIFO_FULL_STATE = 3'b110, LOAD_AFTER_FULL = 3'b111;

reg [2:0] present_state, next_state;

//sequential logic for present state with active low reset and active high soft_reset
always@(posedge clk)
begin 
	if(!rst)
		present_state <= DECODE_ADDRESS;
	else if(soft_reset_0 || soft_reset_1 || soft_reset_2)
		present_state <= DECODE_ADDRESS;
	else
		present_state <= next_state;
end

always@(*) begin
case(present_state)
DECODE_ADDRESS: if((pkt_valid & (data_in[1:0] == 2'b0) & fifo_empty_0) |
				   (pkt_valid & (data_in[1:0] == 2'b01) & fifo_empty_1) |
				   (pkt_valid & (data_in[1:0] == 2'b10) & fifo_empty_2))
				   next_state = LOAD_FIRST_DATA;
				else if((pkt_valid & (data_in[1:0] == 2'b0) & !fifo_empty_0) |
				   (pkt_valid & (data_in[1:0] == 2'b01) & !fifo_empty_1) |
				   (pkt_valid & (data_in[1:0] == 2'b10) & !fifo_empty_2))
				   next_state = WAIT_TILL_EMPTY;
				else
					next_state = DECODE_ADDRESS;
					
WAIT_TILL_EMPTY: if((fifo_empty_0 && (data_in[1:0] == 2'b0)) || (fifo_empty_1 && (data_in[1:0] == 2'b01)) ||
				    (fifo_empty_2 && (data_in[1:0] == 2'b10)))
					next_state = LOAD_FIRST_DATA;
				 else
					next_state = WAIT_TILL_EMPTY;

LOAD_FIRST_DATA: next_state = LOAD_DATA;

LOAD_DATA: if(!fifo_full && !pkt_valid)
			 next_state = LOAD_PARITY;
		   else if(fifo_full)
		     next_state = FIFO_FULL_STATE;
		   else 
		     next_state = LOAD_DATA;
LOAD_PARITY: next_state = CHECK_PARITY_ERROR;

CHECK_PARITY_ERROR: if(fifo_full)
						next_state = FIFO_FULL_STATE;
					else
						next_state = DECODE_ADDRESS;
						
FIFO_FULL_STATE: if(!fifo_full)
					next_state = LOAD_AFTER_FULL;
				 else if(fifo_full)
					next_state = FIFO_FULL_STATE;
					
LOAD_AFTER_FULL: if(!parity_done && low_pkt_valid)
					next_state = LOAD_PARITY;
				 else if(!parity_done && !low_pkt_valid)
					next_state = LOAD_DATA;
				 else if(parity_done)
					next_state = DECODE_ADDRESS;
endcase
end

//Coding style 1 :- Continous assignments for outputs

assign busy = !(present_state == LOAD_DATA || present_state == LOAD_PARITY || present_state == DECODE_ADDRESS);
assign detect_add = (present_state == DECODE_ADDRESS);
assign ld_state = (present_state == LOAD_DATA);
assign laf_state = (present_state == LOAD_AFTER_FULL);
assign full_state = (present_state == FIFO_FULL_STATE);
assign write_enb_reg = (present_state == LOAD_DATA || present_state == LOAD_PARITY || present_state == LOAD_AFTER_FULL);
assign rst_int_reg = (present_state == CHECK_PARITY_ERROR);
assign lfd_state = (present_state == LOAD_FIRST_DATA);


/*
always@(posedge clk) begin
if(!rst || (soft_reset_0 || soft_reset_1 || soft_reset_2)) begin
		busy <= 1'b0;
		detect_add <= 1'b0;
		ld_state <= 1'b0;
		laf_state <= 1'b0;
		full_state <= 1'b0;
		write_enb_reg <= 1'b0;
		rst_int_reg <= 1'b0;
		lfd_state <= 1'b0;
end
else begin
	busy <= 1'b1;
	detect_add <= 1'b0;
		ld_state <= 1'b0;
		laf_state <= 1'b0;
		full_state <= 1'b0;
		write_enb_reg <= 1'b0;
		rst_int_reg <= 1'b0;
		lfd_state <= 1'b0;
	case(present_state)
	DECODE_ADDRESS: detect_add <= 1'b1;
	LOAD_FIRST_DATA: lfd_state <= 1'b1;
	LOAD_DATA: begin 
				busy <= 1'b0;
				ld_state <= 1'b1;
				write_enb_reg <= 1'b1;
			end
	LOAD_PARITY: begin
					busy <= 1'b0;
					write_enb_reg <= 1'b1;
			end
	CHECK_PARITY_ERROR: rst_int_reg <= 1'b1;
	FIFO_FULL_STATE: full_state <= 1'b1;
	LOAD_AFTER_FULL: begin
						write_enb_reg <= 1'b1;
						laf_state <= 1'b1;
					end
	endcase
end
end
*/

endmodule

